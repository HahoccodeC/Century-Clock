module LED7 (
input [3:0] in,
output [6:0] led
);
assign led=(in==0)?7'b0000001: //0
           (in==1)?7'b1001111: //1
			  (in==2)?7'b0010010: //2
			  (in==3)?7'b0000110: //3
			  (in==4)?7'b1001100: //4
			  (in==5)?7'b0100100: //5
			  (in==6)?7'b0100000: //6
			  (in==7)?7'b0001111: //7
			  (in==8)?7'b0000000: //8
			  (in==9)?7'b0000100: //9
			  (in==10)?7'b0001000: //A
			  (in==11)?7'b1100000: //B
			  (in==12)?7'b0110001: //C
			  (in==13)?7'b1000010: //D
			  (in==14)?7'b0110000: //E
			  (in==15)?7'b0111000:7'b0111000; //F
			  
			  
			  
endmodule














